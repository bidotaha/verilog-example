module mulyiplexer_2x1 ( output F,
                         input [1:0] I , S);
wire [1:0] W;
wire Sn;

not (Sn,S);
and (W[0],I[0],Sn);
and (W[1],I[1],S);
or (F,W[1],W[0]);

endmodule 

module multiplexer_2x1_ts();

reg [1:0] I;
reg S;
wire D;

mulyiplexer_2x1 c(D,I,S);

initial
begin

S = 1'b0;
I = 2'b0;

$monitor ("in = %d S = %b out = %b",I,S,D); 

#10 
S = 0; I[0] = 0; I[1] = 1;
#10 
S = 0; I[0] = 1; I[1] = 0;
#10 
S = 1; I[0] = 1; I[1] = 0;
#10 
S = 1; I[0] = 0; I[1] = 1;

end

endmodule  

/////////////////////////////////////////////////////

module mulyiplexer_8x1 ( output F,
                         input [7:0] I , input [2:0] S);
wire [7:0] C;
wire [2:0] Sn;

not (Sn[0],S[0]);
not (Sn[1],S[1]);
not (Sn[2],S[2]);
and (C[0],I[0],Sn[2],Sn[1],Sn[0]);
and (C[1],I[1],Sn[2],Sn[1],S[0]);
and (C[2],I[2],Sn[2],S[1],Sn[0]);
and (C[3],I[3],Sn[2],S[1],S[0]);
and (C[4],I[4],S[2],Sn[1],Sn[0]);
and (C[5],I[5],S[2],Sn[1],S[0]);
and (C[6],I[6],S[2],S[1],Sn[0]);
and (C[7],I[7],S[2],S[1],S[0]);
or (F,C[0],C[1],C[2],C[3],C[4],C[5],C[6],C[7]);

endmodule 


module multiplexer_8x1_ts();

reg [7:0] I;
reg [2:0] S;
wire D;

mulyiplexer_8x1 c(D,I,S);

initial
begin

S = 3'b0;
I = 8'b0;

$monitor ("in = %b S = %b out = %b",I,S,D); 

#10 
S = 3'b000; I[0]=1; I[1]=0; I[2]=0; I[3]=0; I[4]=0; I[5]=0; I[6]=0; I[7]=0;
#10 
S = 3'b001; I[0]=0; I[1]=0; I[2]=0; I[3]=0; I[4]=0; I[5]=0; I[6]=0; I[7]=0;
#10 
S = 3'b010; I[0]=0; I[1]=0; I[2]=1; I[3]=0; I[4]=0; I[5]=0; I[6]=0; I[7]=0;
#10 
S = 3'b011; I[0]=1; I[1]=0; I[2]=0; I[3]=0; I[4]=0; I[5]=0; I[6]=0; I[7]=0;
#10 
S = 3'b100; I[0]=1; I[1]=0; I[2]=0; I[3]=0; I[4]=1; I[5]=0; I[6]=0; I[7]=0;
#10 
S = 3'b101; I[0]=1; I[1]=0; I[2]=0; I[3]=0; I[4]=0; I[5]=0; I[6]=0; I[7]=0;
#10 
S = 3'b110; I[0]=1; I[1]=0; I[2]=0; I[3]=0; I[4]=0; I[5]=0; I[6]=1; I[7]=0;
#10 
S = 3'b111; I[0]=1; I[1]=0; I[2]=0; I[3]=0; I[4]=0; I[5]=0; I[6]=0; I[7]=0;

end

endmodule  

/////////////////////////////////////

module mulyiplexer_16x1 ( output F,
                          input [15:0] I , input [3:0] S);
wire [1:0] W;

mulyiplexer_8x1 C0 (W[0],I[7:0],S[2:0]);
mulyiplexer_8x1 C1 (W[1],I[15:8],S[2:0]);
mulyiplexer_2x1 C3 (F,W,S[3]);

endmodule 

module multiplexer_16x1_ts();

reg [15:0] I;
reg [3:0] S;
wire D;

mulyiplexer_16x1 c(D,I,S);

initial
begin

S = 4'b0;
I = 16'b0;

$monitor ("in = %b S = %b out = %b",I,S,D); 

#10 
S = 4'b0000; I[0]=1; I[1]=0; I[2]=0; I[3]=0; I[4]=0; I[5]=0; I[6]=0; I[7]=0;
#10 
S = 4'b0001; I[0]=0; I[1]=0; I[2]=0; I[3]=0; I[4]=0; I[5]=0; I[6]=0; I[7]=0;
#10 
S = 4'b0010; I[0]=0; I[1]=0; I[2]=1; I[3]=0; I[4]=0; I[5]=0; I[6]=0; I[7]=0;
#10 
S = 4'b0011; I[0]=1; I[1]=0; I[2]=0; I[3]=0; I[4]=0; I[5]=0; I[6]=0; I[7]=0;
#10 
S = 4'b0100; I[0]=1; I[1]=0; I[2]=0; I[3]=0; I[4]=1; I[5]=0; I[6]=0; I[7]=0;
#10 
S = 4'b0101; I[0]=1; I[1]=0; I[2]=0; I[3]=0; I[4]=0; I[5]=0; I[6]=0; I[7]=0;
#10 
S = 4'b0110; I[0]=1; I[1]=0; I[2]=0; I[3]=0; I[4]=0; I[5]=0; I[6]=1; I[7]=0;
#10 
S = 4'b0111; I[0]=1; I[1]=0; I[2]=0; I[3]=0; I[4]=0; I[5]=0; I[6]=0; I[7]=0;
#10 
S = 4'b1000; I[8]=1; I[9]=0; I[10]=0; I[11]=0; I[12]=0; I[13]=0; I[14]=0; I[15]=0;
#10 
S = 4'b1001; I[8]=0; I[9]=1; I[10]=0; I[11]=0; I[12]=0; I[13]=0; I[14]=0; I[15]=0;
#10 
S = 4'b1010; I[8]=0; I[9]=0; I[10]=1; I[11]=0; I[12]=0; I[13]=0; I[14]=0; I[15]=0;
#10 
S = 4'b1011; I[8]=0; I[9]=0; I[10]=0; I[11]=1; I[12]=0; I[13]=0; I[14]=0; I[15]=0;
#10 
S = 4'b1100; I[8]=0; I[9]=0; I[10]=0; I[11]=0; I[12]=1; I[13]=0; I[14]=0; I[15]=0;
#10 
S = 4'b1101; I[8]=0; I[9]=0; I[10]=0; I[11]=0; I[12]=0; I[13]=1; I[14]=0; I[15]=0;
#10 
S = 4'b1110; I[8]=0; I[9]=0; I[10]=0; I[11]=0; I[12]=0; I[13]=0; I[14]=1; I[15]=0;
#10 
S = 4'b1111; I[8]=0; I[9]=0; I[10]=0; I[11]=0; I[12]=0; I[13]=0; I[14]=0; I[15]=1;
end 

endmodule 